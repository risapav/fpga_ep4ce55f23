
---

## 🧰 Voliteľné rozšírenia:

### 1. **MkDocs** – generovanie webovej dokumentácie z Markdownu
- [https://www.mkdocs.org/](https://www.mkdocs.org/)
- Možnosť hostovania cez GitHub Pages

### 2. **Doxygen** (s podporou SystemVerilogu)
- Možné anotovať zdrojové súbory komentármi `///`, `/*! */` a generovať HTML dokumentáciu
- Viac formálne, výhodné pri veľkých projektoch

### 3. **Sphinx + Breathe + Exhale** – ak chceš pokročilejšiu dokumentáciu (vyžaduje viac konfigurácie)

---

## 🧪 Odporúčanie:
- **Začni s Markdownom** v Git repozitári: rýchle, jednoduché, rozšíriteľné.
- Neskôr môžeš dokumentáciu rozšíriť pomocou **MkDocs** alebo **Doxygen**, ak projekt narastie.

---

Ak chceš, môžem ti pripraviť šablónu s úvodným `README.md` a jedným návodom v `docs/`. Chceš?
